// Author: Ciro Fabian Bermudez Marquez
// Name: dec7seg.v
//
// Descrition: 7-Segment Decoder Active high

module top (
  input            clk_i,
  input            rst_i,
  output reg [6:0] seg_o,
  output           dp_o
);


endmodule
