// Author: Ciro Fabian Bermudez Marquez
// Name: rom.v
//
// ROM with all required values A(a , b ) = A(10,21)
module rom #(
   parameter Width = 32
) (
    output [Width-1:0] a_o,
    output [Width-1:0] b_o,
    output [Width-1:0] c_o,
	output [Width-1:0] h_o,
	output [Width-1:0] x0_o,
	output [Width-1:0] y0_o,
	output [Width-1:0] z0_o
);

    assign     a_o = 32'b00000101000000000000000000000000; //   40.0000000000000000000000000
	assign     b_o = 32'b00000011100000000000000000000000; //   28.0000000000000000000000000
	assign     c_o = 32'b00000000011000000000000000000000; //    3.0000000000000000000000000
	assign     h_o = 32'b00000000000000000010100011110101; //    0.0049996376037597656250000
	assign    x0_o = 32'b11111111111111001100110011001101; //   -0.0999999046325683593750000
	assign    y0_o = 32'b00000000000100000000000000000000; //    0.5000000000000000000000000
	assign    z0_o = 32'b11111111111011001100110011001101; //   -0.5999999046325683593750000

endmodule
