// A(7,28)
module rom_coef #(
  parameter  Addr = 6,
  parameter Width = 36
) (
  input       [Addr-1:0] addr_i,
  output reg [Width-1:0] value_o
);
	
	always@(i_i)
		case(i_i)			
			 0: an_o = 36'b111111111010111111101110100001000001; //   -0.00977396208327263593673706054687500 
			 1: an_o = 36'b111111111001010011101001101011011010; //   -0.01307216729037463665008544921875000 
			 2: an_o = 36'b111111110101111001101101000010111100; //   -0.01972339348867535591125488281250000 
			 3: an_o = 36'b111111110011011000011011010001010100; //   -0.02464519953355193138122558593750000 
			 4: an_o = 36'b111111110101101000010110001101000100; //   -0.02025308413431048393249511718750000 
			 5: an_o = 36'b000000000000000000000000000000000000; //    0.00000000000000000000000000000000000 
			 6: an_o = 36'b000000010011011000000101001100111010; //    0.03784427721984684467315673828125000 
			 7: an_o = 36'b000000101101000101110010010100011111; //    0.08806720736902207136154174804687500 
			 8: an_o = 36'b000001000111010100101000011111011101; //    0.13930153439287096261978149414062500 
			 9: an_o = 36'b000001011010111110000110100111010110; //    0.17767649400047957897186279296875000 
			10: an_o = 36'b000001100010010000100011001010010011; //    0.19191129726823419332504272460937500 
			11: an_o = 36'b000001011010111110000110100111010110; //    0.17767649400047957897186279296875000 
			12: an_o = 36'b000001000111010100101000011111011101; //    0.13930153439287096261978149414062500 
			13: an_o = 36'b000000101101000101110010010100011111; //    0.08806720736902207136154174804687500 
			14: an_o = 36'b000000010011011000000101001100111010; //    0.03784427721984684467315673828125000 
			15: an_o = 36'b000000000000000000000000000000000000; //    0.00000000000000000000000000000000000 
			16: an_o = 36'b111111110101101000010110001101000100; //   -0.02025308413431048393249511718750000 
			17: an_o = 36'b111111110011011000011011010001010100; //   -0.02464519953355193138122558593750000 
			18: an_o = 36'b111111110101111001101101000010111100; //   -0.01972339348867535591125488281250000 
			19: an_o = 36'b111111111001010011101001101011011010; //   -0.01307216729037463665008544921875000 
			20: an_o = 36'b111111111010111111101110100001000001; //   -0.00977396208327263593673706054687500 
			default: an_o = 36'b000000000000000000000000000000000000; // 0	 	
			
		endcase
endmodule