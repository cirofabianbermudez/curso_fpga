module rom #(
  parameter n = 32,
	parameter m = 4
)	(
	input		    [m-1:0] addr_i,
	output reg	[n-1:0] angulo_o
	);
	
	always @(addr_i) begin
		case(addr_i)		 
       0 : angulo_o = 32'b00101101000000000000000000000000; //  45.0000000000000000000000000
       1 : angulo_o = 32'b00011010100100001010011100110001; //  26.5650511384010314941406250
       2 : angulo_o = 32'b00001110000010010100011101000000; //  14.0362434387207031250000000
       3 : angulo_o = 32'b00000111001000000000000100010010; //   7.1250163316726684570312500
       4 : angulo_o = 32'b00000011100100111000101010100110; //   3.5763343572616577148437500
       5 : angulo_o = 32'b00000001110010100011011110010100; //   1.7899105548858642578125000
       6 : angulo_o = 32'b00000000111001010010101000011010; //   0.8951736688613891601562500
       7 : angulo_o = 32'b00000000011100101001011011010111; //   0.4476141333580017089843750
       8 : angulo_o = 32'b00000000001110010100101110100101; //   0.2238104939460754394531250
       9 : angulo_o = 32'b00000000000111001010010111011001; //   0.1119056344032287597656250
      10 : angulo_o = 32'b00000000000011100101001011101101; //   0.0559528470039367675781250
      11 : angulo_o = 32'b00000000000001110010100101110110; //   0.0279763936996459960937500
      12 : angulo_o = 32'b00000000000000111001010010111011; //   0.0139881968498229980468750
      13 : angulo_o = 32'b00000000000000011100101001011101; //   0.0069940686225891113281250
      14 : angulo_o = 32'b00000000000000001110010100101110; //   0.0034970045089721679687500
      15 : angulo_o = 32'b00000000000000000111001010010111; //   0.0017485022544860839843750
		  default : angulo_o = 32'b00000000000000000000000000000000; 				
		endcase
  end		
	
endmodule