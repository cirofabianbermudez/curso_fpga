module ajuste (
  input      [59:0] r_i,
  input       [5:0] s_i,
  output reg [17:0] y_o	
); 
	
  always@(r_i, s_i) begin
	case(s_i)
       0 : y_o = r_i[17: 0];
       1 : y_o = r_i[18: 1];
       2 : y_o = r_i[19: 2];
       3 : y_o = r_i[20: 3];
       4 : y_o = r_i[21: 4];
       5 : y_o = r_i[22: 5];
       6 : y_o = r_i[23: 6];
       7 : y_o = r_i[24: 7];
       8 : y_o = r_i[25: 8];
       9 : y_o = r_i[26: 9];
      10 : y_o = r_i[27:10];
      11 : y_o = r_i[28:11];
      12 : y_o = r_i[29:12];
      13 : y_o = r_i[30:13];
      14 : y_o = r_i[31:14];
      15 : y_o = r_i[32:15];
      16 : y_o = r_i[33:16];
      17 : y_o = r_i[34:17];
      18 : y_o = r_i[35:18];
      19 : y_o = r_i[36:19];
      20 : y_o = r_i[37:20];
      21 : y_o = r_i[38:21];
      22 : y_o = r_i[39:22];
      23 : y_o = r_i[40:23];
      24 : y_o = r_i[41:24];
      25 : y_o = r_i[42:25];
      26 : y_o = r_i[43:26];
      27 : y_o = r_i[44:27];
      28 : y_o = r_i[45:28];
      29 : y_o = r_i[46:29];
      30 : y_o = r_i[47:30];
      31 : y_o = r_i[48:31];
      32 : y_o = r_i[49:32];
      33 : y_o = r_i[50:33];
      34 : y_o = r_i[51:34];
      35 : y_o = r_i[52:35];
      36 : y_o = r_i[53:36];
      37 : y_o = r_i[54:37];
      38 : y_o = r_i[55:38];
      39 : y_o = r_i[56:39];
      40 : y_o = r_i[57:40];
      41 : y_o = r_i[58:41];
      42 : y_o = r_i[59:42];
      default: y_o = 0;
    endcase		
  end
  
endmodule